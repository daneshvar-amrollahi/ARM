`include "defines.v"

module cache_controller();
endmodule